`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.01.2026 22:12:38
// Design Name: 
// Module Name: ls_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ls_unit(
    input  [31:0] in,        // Data read from data memory
    input  [31:0] in_s,       // Store data from register file
    input  [31:0] address,    // Effective memory address
    input  [4:0]  lsunit,     // Load/Store control encoding

    output [31:0] out,        // Final load-aligned output
    output [31:0] out_s,      // Store-aligned data
    output [3:0]  strobe      // Byte-enable signals
);

    // =========================================================
    // LSUNIT ENCODING
    // =========================================================
    // lsunit[4]   : Valid load/store instruction
    // lsunit[3]   : 0 = Load, 1 = Store
    // lsunit[2:0] : funct3 field
    //
    // funct3:
    // 000 : LB / SB
    // 001 : LH / SH
    // 010 : LW / SW
    // 100 : LBU
    // 101 : LHU
    // =========================================================

    // =========================================================
    // LOAD DATA ALIGNMENT & SIGN EXTENSION
    // =========================================================
    // Based on address offset and funct3

    assign out = (lsunit[4:3] == 2'b10) ?   // Valid LOAD
                 (
                   // -------------------------------------------------
                   // LB (signed)
                   // -------------------------------------------------
                   (lsunit[2:0] == 3'b000) ?
                        ((address[1:0] == 2'b00) ? {{24{in[7]}},  in[7:0]}   :
                         (address[1:0] == 2'b01) ? {{24{in[15]}}, in[15:8]}  :
                         (address[1:0] == 2'b10) ? {{24{in[23]}}, in[23:16]} :
                                                    {{24{in[31]}}, in[31:24]}) :

                   // -------------------------------------------------
                   // LH (signed)
                   // -------------------------------------------------
                   (lsunit[2:0] == 3'b001) ?
                        ((address[1] == 1'b0) ? {{16{in[15]}}, in[15:0]} :
                                                 {{16{in[31]}}, in[31:16]}) :

                   // -------------------------------------------------
                   // LW
                   // -------------------------------------------------
                   (lsunit[2:0] == 3'b010) ? in :

                   // -------------------------------------------------
                   // LBU (unsigned)
                   // -------------------------------------------------
                   (lsunit[2:0] == 3'b100) ?
                        ((address[1:0] == 2'b00) ? {{24{1'b0}}, in[7:0]}   :
                         (address[1:0] == 2'b01) ? {{24{1'b0}}, in[15:8]}  :
                         (address[1:0] == 2'b10) ? {{24{1'b0}}, in[23:16]} :
                                                    {{24{1'b0}}, in[31:24]}) :

                   // -------------------------------------------------
                   // LHU (unsigned)
                   // -------------------------------------------------
                        ((address[1] == 1'b0) ? {{16{1'b0}}, in[15:0]} :
                                                 {{16{1'b0}}, in[31:16]})
                 )
                 : 32'd0;

    // =========================================================
    // STORE BYTE ENABLE (WSTRB)
    // =========================================================
    // Controls which bytes are written to memory

    assign strobe = (lsunit[4:3] == 2'b11) ?   // Valid STORE
                    (
                        (lsunit[2:0] == 3'b000) ? 4'b0001 :  // SB
                        (lsunit[2:0] == 3'b001) ? 4'b0011 :  // SH
                                                    4'b1111   // SW
                    )
                    : 4'b1111;

    // =========================================================
    // STORE DATA ALIGNMENT
    // =========================================================
    // Aligns register data based on address offset

    assign out_s = (lsunit[4:3] == 2'b11) ?    // Valid STORE
                   (
                       // -------------------------------------------------
                       // SB
                       // -------------------------------------------------
                       (lsunit[2:0] == 3'b000) ?
                            ((address[1:0] == 2'b00) ? in_s :
                             (address[1:0] == 2'b01) ? (in_s << 8)  :
                             (address[1:0] == 2'b10) ? (in_s << 16) :
                                                        (in_s << 24)) :

                       // -------------------------------------------------
                       // SH
                       // -------------------------------------------------
                       (lsunit[2:0] == 3'b001) ?
                            ((address[1] == 1'b0) ? in_s :
                                                     (in_s << 16)) :

                       // -------------------------------------------------
                       // SW
                       // -------------------------------------------------
                       in_s
                   )
                   : in_s;

endmodule
